LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.numeric_std.ALL;
----------------------------------------------------------------------------------
ENTITY MEM IS
    PORT (
        ADDRESS : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
        DATA : OUT STD_LOGIC_VECTOR (5 DOWNTO 0));
END MEM;
----------------------------------------------------------------------------------
ARCHITECTURE Behavioral OF MEM IS
    ----------------------------------------------------------------------------------
    TYPE mem_array IS ARRAY(0 TO 63) OF STD_LOGIC_VECTOR(5 DOWNTO 0);
    CONSTANT ROM : mem_array := (
        --------------TEST Loop (second part of project) ----------------------
        -- 8x6 = 6 times add 8 to 8
        "000011", -- Load R0
        "000000", -- 0
        "000111", -- Load R1
        "000001", -- 1     
        "001011", -- Load R2 (counter)
        "000110", -- 6
        "001111", -- Load R3
        "001000", -- 8
        "010010", -- Add R0, R2 (mem[8])
        "101101", -- Sub R3, R1
        "111011", -- JNZ R3
        "001000", -- 8 (go to mem[8])
        -- "000000", -- HLT (commented this so cpu can continue working)
        --------------reseting registers ----------------------
        "000011", -- Load R0
        "000000", -- 0
        "000100", -- Load R1
        "000000", -- 0
        -- "000000", -- HLT (commented this so cpu can continue working)
        --------------TEST Add (first part of project) ----------------------
        "000011", -- load R0
        "000111", -- 7
        "000111", -- load R1
        "000100", -- 4
        "010001", -- Add R0, R1	
        "000000", -- HLT		  
        "000000",
        "000000",
        "000000",
        "000000",
        "000000",
        "000000",
        "000000",
        "000000",
        "000000",
        "000000",
        "000000",
        "000000",
        "000000",
        "000000",
        "000000",
        "000000",
        "000000",
        "000000",
        "000000",
        "000000",
        "000000",
        "000000",
        "000000",
        "000000",
        "000000",
        "000000",
        "000000",
        "000000",
        "000000",
        "000000",
        "000000",
        "000000",
        "000000",
        "000000",
        "000000",
        "000000",
        "000000",
        "000000",
        "000000",
        "000000",
        "000000",
        "000000"
    );
    ----------------------------------------------------------------------------------
BEGIN
    ----------------------------------------------------------------------------------
    pr : PROCESS (ADDRESS)
    BEGIN
        DATA <= ROM(to_integer(unsigned(ADDRESS(5 DOWNTO 0))));
    END PROCESS; -- pr
    ----------------------------------------------------------------------------------
    ----------------------------------------------------------------------------------
END Behavioral;